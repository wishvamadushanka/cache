module data_mem(
    parameters
) (
    ports
);
    
endmodule